module router ();

endmodule