module 4_stage_processor (
  
);

endmodule